* SPICE3 file created from pfet.ext - technology: sky130A

.option scale=5000u

X0 a_400_0# a_0_n26# a_n60_0# w_n96_n36# sky130_fd_pr__pfet_01v8_lvt w=1000 l=400
